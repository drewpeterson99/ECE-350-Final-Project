module register_64(out, in, clk, clr, en);
    input clk, clr, en;
    input [63:0] in;
    output [63:0] out;

    dffe_ref flop0(out[0], in[0], clk, en, clr);
    dffe_ref flop1(out[1], in[1], clk, en, clr);
    dffe_ref flop2(out[2], in[2], clk, en, clr);
    dffe_ref flop3(out[3], in[3], clk, en, clr);
    dffe_ref flop4(out[4], in[4], clk, en, clr);
    dffe_ref flop5(out[5], in[5], clk, en, clr);
    dffe_ref flop6(out[6], in[6], clk, en, clr);
    dffe_ref flop7(out[7], in[7], clk, en, clr);
    dffe_ref flop8(out[8], in[8], clk, en, clr);
    dffe_ref flop9(out[9], in[9], clk, en, clr);
    dffe_ref flop10(out[10], in[10], clk, en, clr);
    dffe_ref flop11(out[11], in[11], clk, en, clr);
    dffe_ref flop12(out[12], in[12], clk, en, clr);
    dffe_ref flop13(out[13], in[13], clk, en, clr);
    dffe_ref flop14(out[14], in[14], clk, en, clr);
    dffe_ref flop15(out[15], in[15], clk, en, clr);
    dffe_ref flop16(out[16], in[16], clk, en, clr);
    dffe_ref flop17(out[17], in[17], clk, en, clr);
    dffe_ref flop18(out[18], in[18], clk, en, clr);
    dffe_ref flop19(out[19], in[19], clk, en, clr);
    dffe_ref flop20(out[20], in[20], clk, en, clr);
    dffe_ref flop21(out[21], in[21], clk, en, clr);
    dffe_ref flop22(out[22], in[22], clk, en, clr);
    dffe_ref flop23(out[23], in[23], clk, en, clr);
    dffe_ref flop24(out[24], in[24], clk, en, clr);
    dffe_ref flop25(out[25], in[25], clk, en, clr);
    dffe_ref flop26(out[26], in[26], clk, en, clr);
    dffe_ref flop27(out[27], in[27], clk, en, clr);
    dffe_ref flop28(out[28], in[28], clk, en, clr);
    dffe_ref flop29(out[29], in[29], clk, en, clr);
    dffe_ref flop30(out[30], in[30], clk, en, clr);
    dffe_ref flop31(out[31], in[31], clk, en, clr);
    dffe_ref flop32(out[32], in[32], clk, en, clr);
    dffe_ref flop33(out[33], in[33], clk, en, clr);
    dffe_ref flop34(out[34], in[34], clk, en, clr);
    dffe_ref flop35(out[35], in[35], clk, en, clr);
    dffe_ref flop36(out[36], in[36], clk, en, clr);
    dffe_ref flop37(out[37], in[37], clk, en, clr);
    dffe_ref flop38(out[38], in[38], clk, en, clr);
    dffe_ref flop39(out[39], in[39], clk, en, clr);
    dffe_ref flop40(out[40], in[40], clk, en, clr);
    dffe_ref flop41(out[41], in[41], clk, en, clr);
    dffe_ref flop42(out[42], in[42], clk, en, clr);
    dffe_ref flop43(out[43], in[43], clk, en, clr);
    dffe_ref flop44(out[44], in[44], clk, en, clr);
    dffe_ref flop45(out[45], in[45], clk, en, clr);
    dffe_ref flop46(out[46], in[46], clk, en, clr);
    dffe_ref flop47(out[47], in[47], clk, en, clr);
    dffe_ref flop48(out[48], in[48], clk, en, clr);
    dffe_ref flop49(out[49], in[49], clk, en, clr);
    dffe_ref flop50(out[50], in[50], clk, en, clr);
    dffe_ref flop51(out[51], in[51], clk, en, clr);
    dffe_ref flop52(out[52], in[52], clk, en, clr);
    dffe_ref flop53(out[53], in[53], clk, en, clr);
    dffe_ref flop54(out[54], in[54], clk, en, clr);
    dffe_ref flop55(out[55], in[55], clk, en, clr);
    dffe_ref flop56(out[56], in[56], clk, en, clr);
    dffe_ref flop57(out[57], in[57], clk, en, clr);
    dffe_ref flop58(out[58], in[58], clk, en, clr);
    dffe_ref flop59(out[59], in[59], clk, en, clr);
    dffe_ref flop60(out[60], in[60], clk, en, clr);
    dffe_ref flop61(out[61], in[61], clk, en, clr);
    dffe_ref flop62(out[62], in[62], clk, en, clr);
    dffe_ref flop63(out[63], in[63], clk, en, clr);

endmodule